library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity multiplier_eight is
    port(A : in STD_LOGIC_VECTOR(15 downto 0);
         B : in STD_LOGIC_VECTOR(15 downto 0);
         res : out STD_LOGIC_VECTOR(15 downto 0)
     );
end multiplier_eight;

architecture dataflow of multiplier_eight is
    component array_multiplier is
        port(a : in STD_LOGIC_VECTOR(3 downto 0);
             b : in STD_LOGIC_VECTOR(3 downto 0);
             ans : out STD_LOGIC_VECTOR(7 downto 0)
         );
    end component;
    component ripple_sixteen_adder is
    port (A,B:in STD_LOGIC_VECTOR(15 downto 0);
          sum:out STD_LOGIC_VECTOR(15 downto 0);
          cout:out STD_LOGIC;
          command:in STD_LOGIC);
    end component;

    signal s1, s2, s3, s4 : STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";
    signal mid1, mid2 : STD_LOGIC_VECTOR(15 downto 0);
    signal cout1 : STD_LOGIC;
    signal cout2 : STD_LOGIC;
    signal cout3 : STD_LOGIC;
begin
    AM1 : array_multiplier port map(A(3 downto 0), B(3 downto 0), s1(7 downto 0));
    AM2 : array_multiplier port map(A(7 downto 4), B(3 downto 0), s2(11 downto 4));
    AM3 : array_multiplier port map(A(3 downto 0), B(7 downto 4), s3(11 downto 4));
    AM4 : array_multiplier port map(A(7 downto 4), B(7 downto 4), s4(15 downto 8));

    SUM1: ripple_sixteen_adder port map(s1, s2, mid1, cout1, '0');
    SUM2: ripple_sixteen_adder port map(s3, s4, mid2, cout2, '0');
    SUM3: ripple_sixteen_adder port map(mid1, mid2, res,cout3, '0');

end dataflow;
